`ifndef __RGGEN_RAL_PKG_SV__
`define __RGGEN_RAL_PKG_SV__
package rggen_ral_pkg;
  import  uvm_pkg::*;
  `include  "uvm_macros.svh"

  `include  "rggen_ral_macros.svh"
  `include  "rggen_ral_field.svh"
  `include  "rggen_ral_field_rwl_rwe.svh"
  `include  "rggen_ral_reg.svh"
  `include  "rggen_ral_indirect_reg.svh"
  `include  "rggen_ral_map.svh"
  `include  "rggen_ral_block.svh"
endpackage
`endif
