`ifndef __RGEN_RAL_PKG_SV__
`define __RGEN_RAL_PKG_SV__
package rgen_ral_pkg;
  import  uvm_pkg::*;
  `include  "uvm_macros.svh"

  `include  "rgen_ral_macros.svh"
  `include  "rgen_ral_field.svh"
  `include  "rgen_ral_reg.svh"
  `include  "rgen_ral_shadow_reg.svh"
  `include  "rgen_ral_map.svh"
  `include  "rgen_ral_block.svh"
endpackage
`endif
